`timescale 1ns/100ps

module tb_hsv2rgb;
    logic clock = 1'b0;
    logic reset = 1'b1;

    /* Master clock 100MHz (10ns period) */
    always #(10ns/2) clock <= ~clock;

    logic [7:0] h, s, v;
    logic [7:0] r, g, b;
    logic valid, ready;

    hsv2rgb DUT
      (.clock, .reset,
       .h, .s, .v,
       .ready_i(ready),
       .r, .g, .b,
       .valid_o(valid));

    always_ff @ (posedge clock)
      if (valid)
        $display("%d %d %d", r, g, b);

    initial begin
        reset = 1'b1;
        ready = 1'b0;
        repeat(10) @(posedge clock) #1;
        reset = 1'b0;

        @(posedge clock) #1;
        h = 8'd50;
        s = 8'd100;
        v = 8'd150;
        ready = 1'b1;

        @(posedge clock) #1;
        h = 8'dx;
        s = 8'dx;
        v = 8'dx;
        ready = 1'b0;

        @(posedge clock) #1;
        @(posedge clock) #1;
        @(posedge clock) #1;

        @(posedge clock) #1;
        h = 8'd50;
        s = 8'd100;
        v = 8'd150;
        ready = 1'b1;

        @(posedge clock) #1;
        h = 8'd111;
        s = 8'd222;
        v = 8'd33;
        ready = 1'b1;

        @(posedge clock) #1;
        h = 8'd200;
        s = 8'd150;
        v = 8'd50;
        ready = 1'b1;

        @(posedge clock) #1;
        ready = 1'b0;


        repeat(10) @(posedge clock);
        $finish;
    end

    initial begin
        $dumpfile("tb_hsv2rgb.vcd");
        $dumpvars;
    end

endmodule // tb_hsv2rgb
